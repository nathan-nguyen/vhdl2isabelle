architecture PRE of PRE is


begin
end;
  stimulus : process
    begin
      idbits_out <= IDBITS - 1;
    end process stimulus;